module mux2to1(
    input wire a,
    input wire b,
    input wire sel, 
    output wire y
);
    assign y = sel ? b : a; // explicit logic: y = (a & ~sel) | (b & sel);
endmodule